module my_and_gate (
    input a,    // First input
    input b,    // Second input
    output y    // Output
);

    // Bitwise AND operator (&)
    assign y = a & b;

endmodule