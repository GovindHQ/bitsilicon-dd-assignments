module tb_stopwatch;
reg clk =0;
always #10 clk = ~clk;
reg rst_n,start,stop,reset;
wire [7:0] minutes;
wire [5:0] seconds;
wire [1:0] status;

stopwatch_top dut(
    .clk(clk),
    .rst_n(rst_n),
    .start(start),
    .stop(stop),
    .reset(reset),
    .minutes(minutes),
    .seconds(seconds),
    .status(status)
);

initial begin
    rst_n = 0; start = 0; stop = 0; reset = 0;
    #20 rst_n = 1;

    #10 start = 1; #10 start = 0;
    #200;

    stop = 1; #10 stop = 0;
    #50;

    start = 1; #10 start = 0;
    #100;

    reset = 1; #10 reset = 0;
    #50;

    $finish;
end
endmodule
