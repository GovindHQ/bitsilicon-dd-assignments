module my_or_gate (
    input a,
    input b,
    output y
);

    //Bitwise OR operator (|)
    assign y = a | b;

endmodule