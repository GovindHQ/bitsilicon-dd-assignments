module my_xor_gate (
    input a,
    input b,
    output y
);

    //Bitwise XOR operator (^)
    assign y = a ^ b;

endmodule